/* -------- Instruction Decoder --------- */

`default_nettype none
`include "instructions.v"

module Decoder (
    // Inputs
    input wire [31:0] HexCode, // machine code, 8-digit hexdecimal
    // Outputs
    // 1. operands of this instruction
    output wire [4:0] rs, 
    output wire [4:0] rt,
    output wire [4:0] rd, 
    output wire [4:0] shamt, 
    output wire [15:0] imm, 
    output wire [25:0] jaddr,
    // 2. the identity of this instruction
    output wire [`InstrID_WIDTH-1:0] instr_id
);
    // split the bus
    wire [5:0] opcode, funct;
    assign opcode = HexCode[31:26];
    assign rs = HexCode[25:21];
    assign rt = HexCode[20:16];
    assign rd = HexCode[15:11];
    assign shamt = HexCode[10:6];
    assign funct = HexCode[5:0];
    assign imm = HexCode[15:0];
    assign jaddr = HexCode[25:0];

    function [`InstrID_WIDTH-1:0] RType;
        input [5:0] funct;
        begin
            case (funct)
            // Generated By C/C++ Program
            6'h20   :   RType = `ADD      ;
            6'h21   :   RType = `ADDU     ;
            6'h22   :   RType = `SUB      ;
            6'h23   :   RType = `SUBU     ;
            6'h2a   :   RType = `SLT      ;
            6'h2b   :   RType = `SLTU     ;
            6'h24   :   RType = `AND      ;
            6'h25   :   RType = `OR       ;
            6'h26   :   RType = `XOR      ;
            6'h27   :   RType = `NOR      ;
            // Shift Instructions
            6'h0    :   RType = `SLL      ;
            6'h2    :   RType = `SRL      ;
            6'h3    :   RType = `SRA      ;
            6'h4    :   RType = `SLLV     ;
            6'h6    :   RType = `SRLV     ;
            6'h7    :   RType = `SRAV     ;
            // R-Jump Instructions
            6'h8    :   RType = `JR       ;
            6'h9    :   RType = `JALR     ;
            // Default Condition
            default :   RType = 0;
            endcase
        end
    endfunction

    function [`InstrID_WIDTH-1:0] IJType;
        input [5:0] opcode;
        begin
            case (opcode)
            // Generated By C/C++ Program
            6'h08   :   IJType = `ADDI     ;
            6'h09   :   IJType = `ADDIU    ;
            6'h0c   :   IJType = `ANDI     ;
            6'h0d   :   IJType = `ORI      ;
            6'h0e   :   IJType = `XORI     ;
            6'h0f   :   IJType = `LUI      ;
            6'h0a   :   IJType = `SLTI     ;
            6'h0b   :   IJType = `SLTIU    ;
            // Memory Load and Store
            6'h23   :   IJType = `LW       ;
            6'h2b   :   IJType = `SW       ;
            6'h20   :   IJType = `LB       ;
            6'h24   :   IJType = `LBU      ;
            6'h28   :   IJType = `SB       ;
            6'h21   :   IJType = `LH       ;
            6'h25   :   IJType = `LHU      ;
            6'h29   :   IJType = `SH       ;
            // Branch
            6'h04   :   IJType = `BEQ      ;
            6'h05   :   IJType = `BNE      ;
            6'h06   :   IJType = `BLEZ     ;
            6'h07   :   IJType = `BGTZ     ;
            6'h01   :   IJType = `BLTZ     ;
            6'h01   :   IJType = `BGEZ     ;
            // Jump
            6'h02   :   IJType = `J        ;
            6'h03   :   IJType = `JAL      ;
            // Default Condition
            default :   IJType = 0        ;
            endcase
        end
    endfunction
    
    function [`InstrID_WIDTH-1:0] SpecialOp;
        input [4:0] rt;
        begin
            case (rt) 
            5'b00000: SpecialOp = `BLTZ;
            5'b00001: SpecialOp = `BGEZ;
            default: SpecialOp = 0;
            endcase
        end
    endfunction

    assign instr_id = (
        (opcode == 6'b000001) ? (SpecialOp(rt)) : 
        (opcode == 6'b000000) ? (RType(funct)) : 
        (IJType(opcode))
    );

endmodule
