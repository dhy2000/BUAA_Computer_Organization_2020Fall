/* 
 * File Name: mips.v
 * Module Name: mips
 *
 */
`default_nettype none
/* ---------- Includes ---------- */


/* ---------- Main Body ---------- */
module mips (
    input wire clk,
    input wire reset
);
    
endmodule